`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/09/12 16:38:01
// Design Name: 
// Module Name: v_div1k
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module v_div1k(
	input clk,
	output reg div1k
    );
	reg [31:0]divclk_cnt = 0;
	always@(posedge clk) begin
		if()
	end
endmodule
